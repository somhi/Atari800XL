///////////////   GLOBAL DEFINES   ////////////////
	
`define GUEST_TOP atari800_mist_top	// substitute guest_top (lowercase) by guest's Mist top module name		

