library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fce0c287",
    12 => x"86c0c64e",
    13 => x"49fce0c2",
    14 => x"48f0cec2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c3d7",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"d4ff1e4f",
    50 => x"78ffc348",
    51 => x"66c45168",
    52 => x"c888c148",
    53 => x"987058a6",
    54 => x"2687eb05",
    55 => x"1e731e4f",
    56 => x"c34bd4ff",
    57 => x"4a6b7bff",
    58 => x"6b7bffc3",
    59 => x"7232c849",
    60 => x"7bffc3b1",
    61 => x"31c84a6b",
    62 => x"ffc3b271",
    63 => x"c8496b7b",
    64 => x"71b17232",
    65 => x"2687c448",
    66 => x"264c264d",
    67 => x"0e4f264b",
    68 => x"5d5c5b5e",
    69 => x"ff4a710e",
    70 => x"49724cd4",
    71 => x"7199ffc3",
    72 => x"f0cec27c",
    73 => x"87c805bf",
    74 => x"c94866d0",
    75 => x"58a6d430",
    76 => x"d84966d0",
    77 => x"99ffc329",
    78 => x"66d07c71",
    79 => x"c329d049",
    80 => x"7c7199ff",
    81 => x"c84966d0",
    82 => x"99ffc329",
    83 => x"66d07c71",
    84 => x"99ffc349",
    85 => x"49727c71",
    86 => x"ffc329d0",
    87 => x"6c7c7199",
    88 => x"fff0c94b",
    89 => x"abffc34d",
    90 => x"c387d005",
    91 => x"4b6c7cff",
    92 => x"c6028dc1",
    93 => x"abffc387",
    94 => x"7387f002",
    95 => x"87c7fe48",
    96 => x"ff49c01e",
    97 => x"ffc348d4",
    98 => x"c381c178",
    99 => x"04a9b7c8",
   100 => x"4f2687f1",
   101 => x"e71e731e",
   102 => x"dff8c487",
   103 => x"c01ec04b",
   104 => x"f7c1f0ff",
   105 => x"87e7fd49",
   106 => x"a8c186c4",
   107 => x"87eac005",
   108 => x"c348d4ff",
   109 => x"c0c178ff",
   110 => x"c0c0c0c0",
   111 => x"f0e1c01e",
   112 => x"fd49e9c1",
   113 => x"86c487c9",
   114 => x"ca059870",
   115 => x"48d4ff87",
   116 => x"c178ffc3",
   117 => x"fe87cb48",
   118 => x"8bc187e6",
   119 => x"87fdfe05",
   120 => x"e6fc48c0",
   121 => x"1e731e87",
   122 => x"c348d4ff",
   123 => x"4bd378ff",
   124 => x"ffc01ec0",
   125 => x"49c1c1f0",
   126 => x"c487d4fc",
   127 => x"05987086",
   128 => x"d4ff87ca",
   129 => x"78ffc348",
   130 => x"87cb48c1",
   131 => x"c187f1fd",
   132 => x"dbff058b",
   133 => x"fb48c087",
   134 => x"5e0e87f1",
   135 => x"ff0e5c5b",
   136 => x"dbfd4cd4",
   137 => x"1eeac687",
   138 => x"c1f0e1c0",
   139 => x"defb49c8",
   140 => x"c186c487",
   141 => x"87c802a8",
   142 => x"c087eafe",
   143 => x"87e2c148",
   144 => x"7087dafa",
   145 => x"ffffcf49",
   146 => x"a9eac699",
   147 => x"fe87c802",
   148 => x"48c087d3",
   149 => x"c387cbc1",
   150 => x"f1c07cff",
   151 => x"87f4fc4b",
   152 => x"c0029870",
   153 => x"1ec087eb",
   154 => x"c1f0ffc0",
   155 => x"defa49fa",
   156 => x"7086c487",
   157 => x"87d90598",
   158 => x"6c7cffc3",
   159 => x"7cffc349",
   160 => x"c17c7c7c",
   161 => x"c40299c0",
   162 => x"d548c187",
   163 => x"d148c087",
   164 => x"05abc287",
   165 => x"48c087c4",
   166 => x"8bc187c8",
   167 => x"87fdfe05",
   168 => x"e4f948c0",
   169 => x"1e731e87",
   170 => x"48f0cec2",
   171 => x"4bc778c1",
   172 => x"c248d0ff",
   173 => x"87c8fb78",
   174 => x"c348d0ff",
   175 => x"c01ec078",
   176 => x"c0c1d0e5",
   177 => x"87c7f949",
   178 => x"a8c186c4",
   179 => x"4b87c105",
   180 => x"c505abc2",
   181 => x"c048c087",
   182 => x"8bc187f9",
   183 => x"87d0ff05",
   184 => x"c287f7fc",
   185 => x"7058f4ce",
   186 => x"87cd0598",
   187 => x"ffc01ec1",
   188 => x"49d0c1f0",
   189 => x"c487d8f8",
   190 => x"48d4ff86",
   191 => x"c278ffc3",
   192 => x"cec287fe",
   193 => x"d0ff58f8",
   194 => x"ff78c248",
   195 => x"ffc348d4",
   196 => x"f748c178",
   197 => x"ff1e87f5",
   198 => x"d0ff4ad4",
   199 => x"78d1c448",
   200 => x"c17affc3",
   201 => x"87f80589",
   202 => x"731e4f26",
   203 => x"c54b711e",
   204 => x"4adfcdee",
   205 => x"c348d4ff",
   206 => x"486878ff",
   207 => x"02a8fec3",
   208 => x"8ac187c5",
   209 => x"7287ed05",
   210 => x"87c5059a",
   211 => x"eac048c0",
   212 => x"029b7387",
   213 => x"66c887cc",
   214 => x"f549731e",
   215 => x"86c487e7",
   216 => x"66c887c6",
   217 => x"87eefe49",
   218 => x"c348d4ff",
   219 => x"737878ff",
   220 => x"87c5059b",
   221 => x"d048d0ff",
   222 => x"f648c178",
   223 => x"731e87cd",
   224 => x"c04a711e",
   225 => x"48d4ff4b",
   226 => x"ff78ffc3",
   227 => x"c3c448d0",
   228 => x"48d4ff78",
   229 => x"7278ffc3",
   230 => x"f0ffc01e",
   231 => x"f549d1c1",
   232 => x"86c487ed",
   233 => x"cd059870",
   234 => x"1ec0c887",
   235 => x"fd4966cc",
   236 => x"86c487f8",
   237 => x"d0ff4b70",
   238 => x"7378c248",
   239 => x"87cbf548",
   240 => x"5c5b5e0e",
   241 => x"1ec00e5d",
   242 => x"c1f0ffc0",
   243 => x"fef449c9",
   244 => x"c21ed287",
   245 => x"fd49f8ce",
   246 => x"86c887d0",
   247 => x"84c14cc0",
   248 => x"04acb7d2",
   249 => x"cec287f8",
   250 => x"49bf97f8",
   251 => x"c199c0c3",
   252 => x"c005a9c0",
   253 => x"cec287e7",
   254 => x"49bf97ff",
   255 => x"cfc231d0",
   256 => x"4abf97c0",
   257 => x"b17232c8",
   258 => x"97c1cfc2",
   259 => x"71b14abf",
   260 => x"ffffcf4c",
   261 => x"84c19cff",
   262 => x"e7c134ca",
   263 => x"c1cfc287",
   264 => x"c149bf97",
   265 => x"c299c631",
   266 => x"bf97c2cf",
   267 => x"2ab7c74a",
   268 => x"cec2b172",
   269 => x"4abf97fd",
   270 => x"c29dcf4d",
   271 => x"bf97fece",
   272 => x"ca9ac34a",
   273 => x"ffcec232",
   274 => x"c24bbf97",
   275 => x"c2b27333",
   276 => x"bf97c0cf",
   277 => x"9bc0c34b",
   278 => x"732bb7c6",
   279 => x"c181c2b2",
   280 => x"70307148",
   281 => x"7548c149",
   282 => x"724d7030",
   283 => x"7184c14c",
   284 => x"b7c0c894",
   285 => x"87cc06ad",
   286 => x"2db734c1",
   287 => x"adb7c0c8",
   288 => x"87f4ff01",
   289 => x"fef14874",
   290 => x"5b5e0e87",
   291 => x"f80e5d5c",
   292 => x"ded7c286",
   293 => x"c278c048",
   294 => x"c01ed6cf",
   295 => x"87defb49",
   296 => x"987086c4",
   297 => x"c087c505",
   298 => x"87cec948",
   299 => x"7ec14dc0",
   300 => x"bfe9edc0",
   301 => x"ccd0c249",
   302 => x"4bc8714a",
   303 => x"7087ebee",
   304 => x"87c20598",
   305 => x"edc07ec0",
   306 => x"c249bfe5",
   307 => x"714ae8d0",
   308 => x"d5ee4bc8",
   309 => x"05987087",
   310 => x"7ec087c2",
   311 => x"fdc0026e",
   312 => x"dcd6c287",
   313 => x"d7c24dbf",
   314 => x"7ebf9fd4",
   315 => x"ead6c548",
   316 => x"87c705a8",
   317 => x"bfdcd6c2",
   318 => x"6e87ce4d",
   319 => x"d5e9ca48",
   320 => x"87c502a8",
   321 => x"f1c748c0",
   322 => x"d6cfc287",
   323 => x"f949751e",
   324 => x"86c487ec",
   325 => x"c5059870",
   326 => x"c748c087",
   327 => x"edc087dc",
   328 => x"c249bfe5",
   329 => x"714ae8d0",
   330 => x"fdec4bc8",
   331 => x"05987087",
   332 => x"d7c287c8",
   333 => x"78c148de",
   334 => x"edc087da",
   335 => x"c249bfe9",
   336 => x"714accd0",
   337 => x"e1ec4bc8",
   338 => x"02987087",
   339 => x"c087c5c0",
   340 => x"87e6c648",
   341 => x"97d4d7c2",
   342 => x"d5c149bf",
   343 => x"cdc005a9",
   344 => x"d5d7c287",
   345 => x"c249bf97",
   346 => x"c002a9ea",
   347 => x"48c087c5",
   348 => x"c287c7c6",
   349 => x"bf97d6cf",
   350 => x"e9c3487e",
   351 => x"cec002a8",
   352 => x"c3486e87",
   353 => x"c002a8eb",
   354 => x"48c087c5",
   355 => x"c287ebc5",
   356 => x"bf97e1cf",
   357 => x"c0059949",
   358 => x"cfc287cc",
   359 => x"49bf97e2",
   360 => x"c002a9c2",
   361 => x"48c087c5",
   362 => x"c287cfc5",
   363 => x"bf97e3cf",
   364 => x"dad7c248",
   365 => x"484c7058",
   366 => x"d7c288c1",
   367 => x"cfc258de",
   368 => x"49bf97e4",
   369 => x"cfc28175",
   370 => x"4abf97e5",
   371 => x"a17232c8",
   372 => x"ebdbc27e",
   373 => x"c2786e48",
   374 => x"bf97e6cf",
   375 => x"58a6c848",
   376 => x"bfded7c2",
   377 => x"87d4c202",
   378 => x"bfe5edc0",
   379 => x"e8d0c249",
   380 => x"4bc8714a",
   381 => x"7087f3e9",
   382 => x"c5c00298",
   383 => x"c348c087",
   384 => x"d7c287f8",
   385 => x"c24cbfd6",
   386 => x"c25cffdb",
   387 => x"bf97fbcf",
   388 => x"c231c849",
   389 => x"bf97facf",
   390 => x"c249a14a",
   391 => x"bf97fccf",
   392 => x"7232d04a",
   393 => x"cfc249a1",
   394 => x"4abf97fd",
   395 => x"a17232d8",
   396 => x"9166c449",
   397 => x"bfebdbc2",
   398 => x"f3dbc281",
   399 => x"c3d0c259",
   400 => x"c84abf97",
   401 => x"c2d0c232",
   402 => x"a24bbf97",
   403 => x"c4d0c24a",
   404 => x"d04bbf97",
   405 => x"4aa27333",
   406 => x"97c5d0c2",
   407 => x"9bcf4bbf",
   408 => x"a27333d8",
   409 => x"f7dbc24a",
   410 => x"f3dbc25a",
   411 => x"8ac24abf",
   412 => x"dbc29274",
   413 => x"a17248f7",
   414 => x"87cac178",
   415 => x"97e8cfc2",
   416 => x"31c849bf",
   417 => x"97e7cfc2",
   418 => x"49a14abf",
   419 => x"59e6d7c2",
   420 => x"bfe2d7c2",
   421 => x"c731c549",
   422 => x"29c981ff",
   423 => x"59ffdbc2",
   424 => x"97edcfc2",
   425 => x"32c84abf",
   426 => x"97eccfc2",
   427 => x"4aa24bbf",
   428 => x"6e9266c4",
   429 => x"fbdbc282",
   430 => x"f3dbc25a",
   431 => x"c278c048",
   432 => x"7248efdb",
   433 => x"dbc278a1",
   434 => x"dbc248ff",
   435 => x"c278bff3",
   436 => x"c248c3dc",
   437 => x"78bff7db",
   438 => x"bfded7c2",
   439 => x"87c9c002",
   440 => x"30c44874",
   441 => x"c9c07e70",
   442 => x"fbdbc287",
   443 => x"30c448bf",
   444 => x"d7c27e70",
   445 => x"786e48e2",
   446 => x"8ef848c1",
   447 => x"4c264d26",
   448 => x"4f264b26",
   449 => x"5c5b5e0e",
   450 => x"4a710e5d",
   451 => x"bfded7c2",
   452 => x"7287cb02",
   453 => x"722bc74b",
   454 => x"9cffc14c",
   455 => x"4b7287c9",
   456 => x"4c722bc8",
   457 => x"c29cffc3",
   458 => x"83bfebdb",
   459 => x"bfe1edc0",
   460 => x"87d902ab",
   461 => x"5be5edc0",
   462 => x"1ed6cfc2",
   463 => x"fdf04973",
   464 => x"7086c487",
   465 => x"87c50598",
   466 => x"e6c048c0",
   467 => x"ded7c287",
   468 => x"87d202bf",
   469 => x"91c44974",
   470 => x"81d6cfc2",
   471 => x"ffcf4d69",
   472 => x"9dffffff",
   473 => x"497487cb",
   474 => x"cfc291c2",
   475 => x"699f81d6",
   476 => x"fe48754d",
   477 => x"5e0e87c6",
   478 => x"0e5d5c5b",
   479 => x"c04d711e",
   480 => x"c849c11e",
   481 => x"86c487c4",
   482 => x"029c4c70",
   483 => x"c287c0c1",
   484 => x"754ae6d7",
   485 => x"87f7e249",
   486 => x"c0029870",
   487 => x"4a7487f1",
   488 => x"4bcb4975",
   489 => x"7087dde3",
   490 => x"e2c00298",
   491 => x"741ec087",
   492 => x"87c7029c",
   493 => x"c048a6c4",
   494 => x"c487c578",
   495 => x"78c148a6",
   496 => x"c74966c4",
   497 => x"86c487c4",
   498 => x"059c4c70",
   499 => x"7487c0ff",
   500 => x"e7fc2648",
   501 => x"5b5e0e87",
   502 => x"1e0e5d5c",
   503 => x"059b4b71",
   504 => x"48c087c5",
   505 => x"c887e5c1",
   506 => x"7dc04da3",
   507 => x"c70266d4",
   508 => x"9766d487",
   509 => x"87c505bf",
   510 => x"cfc148c0",
   511 => x"4966d487",
   512 => x"7087f3fd",
   513 => x"c1029c4c",
   514 => x"a4dc87c0",
   515 => x"da7d6949",
   516 => x"a3c449a4",
   517 => x"7a699f4a",
   518 => x"bfded7c2",
   519 => x"d487d202",
   520 => x"699f49a4",
   521 => x"ffffc049",
   522 => x"d0487199",
   523 => x"c27e7030",
   524 => x"6e7ec087",
   525 => x"806a4849",
   526 => x"7bc07a70",
   527 => x"6a49a3cc",
   528 => x"49a3d079",
   529 => x"487479c0",
   530 => x"48c087c2",
   531 => x"87ecfa26",
   532 => x"5c5b5e0e",
   533 => x"4c710e5d",
   534 => x"48e1edc0",
   535 => x"9c7478ff",
   536 => x"87cac102",
   537 => x"6949a4c8",
   538 => x"87c2c102",
   539 => x"6c4a66d0",
   540 => x"a6d48249",
   541 => x"4d66d05a",
   542 => x"dad7c2b9",
   543 => x"baff4abf",
   544 => x"99719972",
   545 => x"87e4c002",
   546 => x"6b4ba4c4",
   547 => x"87f4f949",
   548 => x"d7c27b70",
   549 => x"6c49bfd6",
   550 => x"757c7181",
   551 => x"dad7c2b9",
   552 => x"baff4abf",
   553 => x"99719972",
   554 => x"87dcff05",
   555 => x"cbf97c75",
   556 => x"1e731e87",
   557 => x"029b4b71",
   558 => x"a3c887c7",
   559 => x"c5056949",
   560 => x"c048c087",
   561 => x"dbc287eb",
   562 => x"c44abfef",
   563 => x"496949a3",
   564 => x"d7c289c2",
   565 => x"7191bfd6",
   566 => x"d7c24aa2",
   567 => x"6b49bfda",
   568 => x"4aa27199",
   569 => x"721e66c8",
   570 => x"87d2ea49",
   571 => x"497086c4",
   572 => x"87ccf848",
   573 => x"711e731e",
   574 => x"c0029b4b",
   575 => x"dcc287e4",
   576 => x"4a735bc3",
   577 => x"d7c28ac2",
   578 => x"9249bfd6",
   579 => x"bfefdbc2",
   580 => x"c2807248",
   581 => x"7158c7dc",
   582 => x"c230c448",
   583 => x"c058e6d7",
   584 => x"dbc287ed",
   585 => x"dbc248ff",
   586 => x"c278bff3",
   587 => x"c248c3dc",
   588 => x"78bff7db",
   589 => x"bfded7c2",
   590 => x"c287c902",
   591 => x"49bfd6d7",
   592 => x"87c731c4",
   593 => x"bffbdbc2",
   594 => x"c231c449",
   595 => x"f659e6d7",
   596 => x"5e0e87ee",
   597 => x"710e5c5b",
   598 => x"724bc04a",
   599 => x"e1c0029a",
   600 => x"49a2da87",
   601 => x"c24b699f",
   602 => x"02bfded7",
   603 => x"a2d487cf",
   604 => x"49699f49",
   605 => x"ffffc04c",
   606 => x"c234d09c",
   607 => x"744cc087",
   608 => x"4973b349",
   609 => x"f587edfd",
   610 => x"5e0e87f4",
   611 => x"0e5d5c5b",
   612 => x"4a7186f4",
   613 => x"9a727ec0",
   614 => x"c287d802",
   615 => x"c048d2cf",
   616 => x"cacfc278",
   617 => x"c3dcc248",
   618 => x"cfc278bf",
   619 => x"dbc248ce",
   620 => x"c278bfff",
   621 => x"c048f3d7",
   622 => x"e2d7c250",
   623 => x"cfc249bf",
   624 => x"714abfd2",
   625 => x"ffc303aa",
   626 => x"cf497287",
   627 => x"e0c00599",
   628 => x"d6cfc287",
   629 => x"cacfc21e",
   630 => x"cfc249bf",
   631 => x"a1c148ca",
   632 => x"d9e67178",
   633 => x"c086c487",
   634 => x"c248dded",
   635 => x"cc78d6cf",
   636 => x"ddedc087",
   637 => x"e0c048bf",
   638 => x"e1edc080",
   639 => x"d2cfc258",
   640 => x"80c148bf",
   641 => x"58d6cfc2",
   642 => x"000b5d27",
   643 => x"bf97bf00",
   644 => x"c2029d4d",
   645 => x"e5c387e2",
   646 => x"dbc202ad",
   647 => x"ddedc087",
   648 => x"a3cb4bbf",
   649 => x"cf4c1149",
   650 => x"d2c105ac",
   651 => x"df497587",
   652 => x"cd89c199",
   653 => x"e6d7c291",
   654 => x"4aa3c181",
   655 => x"a3c35112",
   656 => x"c551124a",
   657 => x"51124aa3",
   658 => x"124aa3c7",
   659 => x"4aa3c951",
   660 => x"a3ce5112",
   661 => x"d051124a",
   662 => x"51124aa3",
   663 => x"124aa3d2",
   664 => x"4aa3d451",
   665 => x"a3d65112",
   666 => x"d851124a",
   667 => x"51124aa3",
   668 => x"124aa3dc",
   669 => x"4aa3de51",
   670 => x"7ec15112",
   671 => x"7487f9c0",
   672 => x"0599c849",
   673 => x"7487eac0",
   674 => x"0599d049",
   675 => x"66dc87d0",
   676 => x"87cac002",
   677 => x"66dc4973",
   678 => x"0298700f",
   679 => x"056e87d3",
   680 => x"c287c6c0",
   681 => x"c048e6d7",
   682 => x"ddedc050",
   683 => x"e7c248bf",
   684 => x"f3d7c287",
   685 => x"7e50c048",
   686 => x"bfe2d7c2",
   687 => x"d2cfc249",
   688 => x"aa714abf",
   689 => x"87c1fc04",
   690 => x"bfc3dcc2",
   691 => x"87c8c005",
   692 => x"bfded7c2",
   693 => x"87fec102",
   694 => x"48e1edc0",
   695 => x"cfc278ff",
   696 => x"f049bfce",
   697 => x"497087de",
   698 => x"59d2cfc2",
   699 => x"c248a6c4",
   700 => x"78bfcecf",
   701 => x"bfded7c2",
   702 => x"87d8c002",
   703 => x"cf4966c4",
   704 => x"f8ffffff",
   705 => x"c002a999",
   706 => x"4dc087c5",
   707 => x"c187e1c0",
   708 => x"87dcc04d",
   709 => x"cf4966c4",
   710 => x"a999f8ff",
   711 => x"87c8c002",
   712 => x"c048a6c8",
   713 => x"87c5c078",
   714 => x"c148a6c8",
   715 => x"4d66c878",
   716 => x"c0059d75",
   717 => x"66c487e0",
   718 => x"c289c249",
   719 => x"4abfd6d7",
   720 => x"efdbc291",
   721 => x"cfc24abf",
   722 => x"a17248ca",
   723 => x"d2cfc278",
   724 => x"f978c048",
   725 => x"48c087e3",
   726 => x"dfee8ef4",
   727 => x"00000087",
   728 => x"ffffff00",
   729 => x"000b6dff",
   730 => x"000b7600",
   731 => x"54414600",
   732 => x"20203233",
   733 => x"41460020",
   734 => x"20363154",
   735 => x"1e002020",
   736 => x"c348d4ff",
   737 => x"486878ff",
   738 => x"ff1e4f26",
   739 => x"ffc348d4",
   740 => x"48d0ff78",
   741 => x"ff78e1c8",
   742 => x"78d448d4",
   743 => x"48c7dcc2",
   744 => x"50bfd4ff",
   745 => x"ff1e4f26",
   746 => x"e0c048d0",
   747 => x"1e4f2678",
   748 => x"7087ccff",
   749 => x"c6029949",
   750 => x"a9fbc087",
   751 => x"7187f105",
   752 => x"0e4f2648",
   753 => x"0e5c5b5e",
   754 => x"4cc04b71",
   755 => x"7087f0fe",
   756 => x"c0029949",
   757 => x"ecc087f9",
   758 => x"f2c002a9",
   759 => x"a9fbc087",
   760 => x"87ebc002",
   761 => x"acb766cc",
   762 => x"d087c703",
   763 => x"87c20266",
   764 => x"99715371",
   765 => x"c187c202",
   766 => x"87c3fe84",
   767 => x"02994970",
   768 => x"ecc087cd",
   769 => x"87c702a9",
   770 => x"05a9fbc0",
   771 => x"d087d5ff",
   772 => x"87c30266",
   773 => x"c07b97c0",
   774 => x"c405a9ec",
   775 => x"c54a7487",
   776 => x"c04a7487",
   777 => x"48728a0a",
   778 => x"4d2687c2",
   779 => x"4b264c26",
   780 => x"fd1e4f26",
   781 => x"497087c9",
   782 => x"a9b7f0c0",
   783 => x"c087ca04",
   784 => x"01a9b7f9",
   785 => x"f0c087c3",
   786 => x"b7c1c189",
   787 => x"87ca04a9",
   788 => x"a9b7dac1",
   789 => x"c087c301",
   790 => x"487189f7",
   791 => x"5e0e4f26",
   792 => x"710e5c5b",
   793 => x"4cd4ff4a",
   794 => x"eac04972",
   795 => x"9b4b7087",
   796 => x"c187c202",
   797 => x"48d0ff8b",
   798 => x"c178c5c8",
   799 => x"49737cd5",
   800 => x"cdc231c6",
   801 => x"4abf97db",
   802 => x"70b07148",
   803 => x"48d0ff7c",
   804 => x"487378c4",
   805 => x"0e87d5fe",
   806 => x"5d5c5b5e",
   807 => x"7186f80e",
   808 => x"fb7ec04c",
   809 => x"4bc087e4",
   810 => x"97c4f5c0",
   811 => x"a9c049bf",
   812 => x"fb87cf04",
   813 => x"83c187f9",
   814 => x"97c4f5c0",
   815 => x"06ab49bf",
   816 => x"f5c087f1",
   817 => x"02bf97c4",
   818 => x"f2fa87cf",
   819 => x"99497087",
   820 => x"c087c602",
   821 => x"f105a9ec",
   822 => x"fa4bc087",
   823 => x"4d7087e1",
   824 => x"c887dcfa",
   825 => x"d6fa58a6",
   826 => x"c14a7087",
   827 => x"49a4c883",
   828 => x"ad496997",
   829 => x"c087c702",
   830 => x"c005adff",
   831 => x"a4c987e7",
   832 => x"49699749",
   833 => x"02a966c4",
   834 => x"c04887c7",
   835 => x"d405a8ff",
   836 => x"49a4ca87",
   837 => x"aa496997",
   838 => x"c087c602",
   839 => x"c405aaff",
   840 => x"d07ec187",
   841 => x"adecc087",
   842 => x"c087c602",
   843 => x"c405adfb",
   844 => x"c14bc087",
   845 => x"fe026e7e",
   846 => x"e9f987e1",
   847 => x"f8487387",
   848 => x"87e6fb8e",
   849 => x"5b5e0e00",
   850 => x"1e0e5d5c",
   851 => x"4cc04b71",
   852 => x"c004ab4d",
   853 => x"f2c087e8",
   854 => x"9d751ed7",
   855 => x"c087c402",
   856 => x"c187c24a",
   857 => x"f049724a",
   858 => x"86c487e0",
   859 => x"84c17e70",
   860 => x"87c2056e",
   861 => x"85c14c73",
   862 => x"ff06ac73",
   863 => x"486e87d8",
   864 => x"264d2626",
   865 => x"264b264c",
   866 => x"5b5e0e4f",
   867 => x"1e0e5d5c",
   868 => x"de494c71",
   869 => x"e1dcc291",
   870 => x"9785714d",
   871 => x"ddc1026d",
   872 => x"ccdcc287",
   873 => x"82744abf",
   874 => x"d8fe4972",
   875 => x"6e7e7087",
   876 => x"87f3c002",
   877 => x"4bd4dcc2",
   878 => x"49cb4a6e",
   879 => x"87e8cbff",
   880 => x"93cb4b74",
   881 => x"83f2d8c1",
   882 => x"f8c083c4",
   883 => x"49747bc2",
   884 => x"87e9c2c1",
   885 => x"dcc27b75",
   886 => x"49bf97e0",
   887 => x"d4dcc21e",
   888 => x"e7d5c149",
   889 => x"7486c487",
   890 => x"d0c2c149",
   891 => x"c149c087",
   892 => x"c287efc3",
   893 => x"c048c8dc",
   894 => x"dd49c178",
   895 => x"fd2687cb",
   896 => x"6f4c87ff",
   897 => x"6e696461",
   898 => x"2e2e2e67",
   899 => x"5b5e0e00",
   900 => x"4b710e5c",
   901 => x"ccdcc24a",
   902 => x"497282bf",
   903 => x"7087e6fc",
   904 => x"c4029c4c",
   905 => x"e9ec4987",
   906 => x"ccdcc287",
   907 => x"c178c048",
   908 => x"87d5dc49",
   909 => x"0e87ccfd",
   910 => x"5d5c5b5e",
   911 => x"c286f40e",
   912 => x"c04dd6cf",
   913 => x"48a6c44c",
   914 => x"dcc278c0",
   915 => x"c049bfcc",
   916 => x"c1c106a9",
   917 => x"d6cfc287",
   918 => x"c0029848",
   919 => x"f2c087f8",
   920 => x"66c81ed7",
   921 => x"c487c702",
   922 => x"78c048a6",
   923 => x"a6c487c5",
   924 => x"c478c148",
   925 => x"d1ec4966",
   926 => x"7086c487",
   927 => x"c484c14d",
   928 => x"80c14866",
   929 => x"c258a6c8",
   930 => x"49bfccdc",
   931 => x"87c603ac",
   932 => x"ff059d75",
   933 => x"4cc087c8",
   934 => x"c3029d75",
   935 => x"f2c087e0",
   936 => x"66c81ed7",
   937 => x"cc87c702",
   938 => x"78c048a6",
   939 => x"a6cc87c5",
   940 => x"cc78c148",
   941 => x"d1eb4966",
   942 => x"7086c487",
   943 => x"c2026e7e",
   944 => x"496e87e9",
   945 => x"699781cb",
   946 => x"0299d049",
   947 => x"c087d6c1",
   948 => x"744acdf8",
   949 => x"c191cb49",
   950 => x"7281f2d8",
   951 => x"c381c879",
   952 => x"497451ff",
   953 => x"dcc291de",
   954 => x"85714de1",
   955 => x"7d97c1c2",
   956 => x"c049a5c1",
   957 => x"d7c251e0",
   958 => x"02bf97e6",
   959 => x"84c187d2",
   960 => x"c24ba5c2",
   961 => x"db4ae6d7",
   962 => x"dbc6ff49",
   963 => x"87dbc187",
   964 => x"c049a5cd",
   965 => x"c284c151",
   966 => x"4a6e4ba5",
   967 => x"c6ff49cb",
   968 => x"c6c187c6",
   969 => x"c9f6c087",
   970 => x"cb49744a",
   971 => x"f2d8c191",
   972 => x"c2797281",
   973 => x"bf97e6d7",
   974 => x"7487d802",
   975 => x"c191de49",
   976 => x"e1dcc284",
   977 => x"c283714b",
   978 => x"dd4ae6d7",
   979 => x"d7c5ff49",
   980 => x"7487d887",
   981 => x"c293de4b",
   982 => x"cb83e1dc",
   983 => x"51c049a3",
   984 => x"6e7384c1",
   985 => x"ff49cb4a",
   986 => x"c487fdc4",
   987 => x"80c14866",
   988 => x"c758a6c8",
   989 => x"c5c003ac",
   990 => x"fc056e87",
   991 => x"487487e0",
   992 => x"fcf78ef4",
   993 => x"1e731e87",
   994 => x"cb494b71",
   995 => x"f2d8c191",
   996 => x"4aa1c881",
   997 => x"48dbcdc2",
   998 => x"a1c95012",
   999 => x"c4f5c04a",
  1000 => x"ca501248",
  1001 => x"e0dcc281",
  1002 => x"c2501148",
  1003 => x"bf97e0dc",
  1004 => x"49c01e49",
  1005 => x"87d4cec1",
  1006 => x"48c8dcc2",
  1007 => x"49c178de",
  1008 => x"2687c6d6",
  1009 => x"1e87fef6",
  1010 => x"cb494a71",
  1011 => x"f2d8c191",
  1012 => x"1181c881",
  1013 => x"ccdcc248",
  1014 => x"ccdcc258",
  1015 => x"c178c048",
  1016 => x"87e5d549",
  1017 => x"c01e4f26",
  1018 => x"f5fbc049",
  1019 => x"1e4f2687",
  1020 => x"d2029971",
  1021 => x"c7dac187",
  1022 => x"f750c048",
  1023 => x"c7ffc080",
  1024 => x"ebd8c140",
  1025 => x"c187ce78",
  1026 => x"c148c3da",
  1027 => x"fc78e4d8",
  1028 => x"e6ffc080",
  1029 => x"0e4f2678",
  1030 => x"0e5c5b5e",
  1031 => x"cb4a4c71",
  1032 => x"f2d8c192",
  1033 => x"49a2c882",
  1034 => x"974ba2c9",
  1035 => x"971e4b6b",
  1036 => x"ca1e4969",
  1037 => x"c0491282",
  1038 => x"c087f0e6",
  1039 => x"87c9d449",
  1040 => x"f8c04974",
  1041 => x"8ef887f7",
  1042 => x"1e87f8f4",
  1043 => x"4b711e73",
  1044 => x"87c3ff49",
  1045 => x"fefe4973",
  1046 => x"87e9f487",
  1047 => x"711e731e",
  1048 => x"4aa3c64b",
  1049 => x"c187db02",
  1050 => x"87d6028a",
  1051 => x"dac1028a",
  1052 => x"c0028a87",
  1053 => x"028a87fc",
  1054 => x"8a87e1c0",
  1055 => x"c187cb02",
  1056 => x"49c787db",
  1057 => x"c187c0fd",
  1058 => x"dcc287de",
  1059 => x"c102bfcc",
  1060 => x"c14887cb",
  1061 => x"d0dcc288",
  1062 => x"87c1c158",
  1063 => x"bfd0dcc2",
  1064 => x"87f9c002",
  1065 => x"bfccdcc2",
  1066 => x"c280c148",
  1067 => x"c058d0dc",
  1068 => x"dcc287eb",
  1069 => x"c649bfcc",
  1070 => x"d0dcc289",
  1071 => x"a9b7c059",
  1072 => x"c287da03",
  1073 => x"c048ccdc",
  1074 => x"c287d278",
  1075 => x"02bfd0dc",
  1076 => x"dcc287cb",
  1077 => x"c648bfcc",
  1078 => x"d0dcc280",
  1079 => x"d149c058",
  1080 => x"497387e7",
  1081 => x"87d5f6c0",
  1082 => x"0e87daf2",
  1083 => x"0e5c5b5e",
  1084 => x"66cc4c71",
  1085 => x"cb4b741e",
  1086 => x"f2d8c193",
  1087 => x"4aa3c483",
  1088 => x"fefe496a",
  1089 => x"fec087f2",
  1090 => x"a3c87bc5",
  1091 => x"5166d449",
  1092 => x"d849a3c9",
  1093 => x"a3ca5166",
  1094 => x"5166dc49",
  1095 => x"87e3f126",
  1096 => x"5c5b5e0e",
  1097 => x"d0ff0e5d",
  1098 => x"59a6d886",
  1099 => x"c048a6c4",
  1100 => x"c180c478",
  1101 => x"c47866c4",
  1102 => x"c478c180",
  1103 => x"c278c180",
  1104 => x"c148d0dc",
  1105 => x"c8dcc278",
  1106 => x"a8de48bf",
  1107 => x"f387cb05",
  1108 => x"497087e5",
  1109 => x"ce59a6c8",
  1110 => x"ede887f8",
  1111 => x"87cfe987",
  1112 => x"7087dce8",
  1113 => x"acfbc04c",
  1114 => x"87d0c102",
  1115 => x"c10566d4",
  1116 => x"1ec087c2",
  1117 => x"c11ec11e",
  1118 => x"c01ee5da",
  1119 => x"87ebfd49",
  1120 => x"4a66d0c1",
  1121 => x"496a82c4",
  1122 => x"517481c7",
  1123 => x"1ed81ec1",
  1124 => x"81c8496a",
  1125 => x"d887ece8",
  1126 => x"66c4c186",
  1127 => x"01a8c048",
  1128 => x"a6c487c7",
  1129 => x"ce78c148",
  1130 => x"66c4c187",
  1131 => x"cc88c148",
  1132 => x"87c358a6",
  1133 => x"cc87f8e7",
  1134 => x"78c248a6",
  1135 => x"cd029c74",
  1136 => x"66c487cc",
  1137 => x"66c8c148",
  1138 => x"c1cd03a8",
  1139 => x"48a6d887",
  1140 => x"eae678c0",
  1141 => x"c14c7087",
  1142 => x"c205acd0",
  1143 => x"66d887d6",
  1144 => x"87cee97e",
  1145 => x"a6dc4970",
  1146 => x"87d3e659",
  1147 => x"ecc04c70",
  1148 => x"eac105ac",
  1149 => x"4966c487",
  1150 => x"c0c191cb",
  1151 => x"a1c48166",
  1152 => x"c84d6a4a",
  1153 => x"66d84aa1",
  1154 => x"c7ffc052",
  1155 => x"87efe579",
  1156 => x"029c4c70",
  1157 => x"fbc087d8",
  1158 => x"87d202ac",
  1159 => x"dee55574",
  1160 => x"9c4c7087",
  1161 => x"c087c702",
  1162 => x"ff05acfb",
  1163 => x"e0c087ee",
  1164 => x"55c1c255",
  1165 => x"d47d97c0",
  1166 => x"a96e4966",
  1167 => x"c487db05",
  1168 => x"66c84866",
  1169 => x"87ca04a8",
  1170 => x"c14866c4",
  1171 => x"58a6c880",
  1172 => x"66c887c8",
  1173 => x"cc88c148",
  1174 => x"e2e458a6",
  1175 => x"c14c7087",
  1176 => x"c805acd0",
  1177 => x"4866d087",
  1178 => x"a6d480c1",
  1179 => x"acd0c158",
  1180 => x"87eafd02",
  1181 => x"d448a6dc",
  1182 => x"66d87866",
  1183 => x"a866dc48",
  1184 => x"87dcc905",
  1185 => x"48a6e0c0",
  1186 => x"c478f0c0",
  1187 => x"7866cc80",
  1188 => x"78c080c4",
  1189 => x"c048747e",
  1190 => x"f0c088fb",
  1191 => x"987058a6",
  1192 => x"87d7c802",
  1193 => x"c088cb48",
  1194 => x"7058a6f0",
  1195 => x"e9c00298",
  1196 => x"88c94887",
  1197 => x"58a6f0c0",
  1198 => x"c3029870",
  1199 => x"c44887e1",
  1200 => x"a6f0c088",
  1201 => x"02987058",
  1202 => x"c14887d6",
  1203 => x"a6f0c088",
  1204 => x"02987058",
  1205 => x"c787c8c3",
  1206 => x"e0c087db",
  1207 => x"78c048a6",
  1208 => x"c14866cc",
  1209 => x"58a6d080",
  1210 => x"7087d4e2",
  1211 => x"acecc04c",
  1212 => x"c087d502",
  1213 => x"c60266e0",
  1214 => x"a6e4c087",
  1215 => x"7487c95c",
  1216 => x"88f0c048",
  1217 => x"58a6e8c0",
  1218 => x"02acecc0",
  1219 => x"eee187cc",
  1220 => x"c04c7087",
  1221 => x"ff05acec",
  1222 => x"e0c087f4",
  1223 => x"66d41e66",
  1224 => x"ecc01e49",
  1225 => x"dac11e66",
  1226 => x"66d41ee5",
  1227 => x"87fbf649",
  1228 => x"1eca1ec0",
  1229 => x"cb4966dc",
  1230 => x"66d8c191",
  1231 => x"48a6d881",
  1232 => x"d878a1c4",
  1233 => x"e149bf66",
  1234 => x"86d887f9",
  1235 => x"06a8b7c0",
  1236 => x"c187c7c1",
  1237 => x"c81ede1e",
  1238 => x"e149bf66",
  1239 => x"86c887e5",
  1240 => x"c0484970",
  1241 => x"e4c08808",
  1242 => x"b7c058a6",
  1243 => x"e9c006a8",
  1244 => x"66e0c087",
  1245 => x"a8b7dd48",
  1246 => x"6e87df03",
  1247 => x"e0c049bf",
  1248 => x"e0c08166",
  1249 => x"c1496651",
  1250 => x"81bf6e81",
  1251 => x"c051c1c2",
  1252 => x"c24966e0",
  1253 => x"81bf6e81",
  1254 => x"7ec151c0",
  1255 => x"e287dcc4",
  1256 => x"e4c087d0",
  1257 => x"c9e258a6",
  1258 => x"a6e8c087",
  1259 => x"a8ecc058",
  1260 => x"87cbc005",
  1261 => x"48a6e4c0",
  1262 => x"7866e0c0",
  1263 => x"ff87c4c0",
  1264 => x"c487fcde",
  1265 => x"91cb4966",
  1266 => x"4866c0c1",
  1267 => x"7e708071",
  1268 => x"82c84a6e",
  1269 => x"81ca496e",
  1270 => x"5166e0c0",
  1271 => x"4966e4c0",
  1272 => x"e0c081c1",
  1273 => x"48c18966",
  1274 => x"49703071",
  1275 => x"977189c1",
  1276 => x"fddfc27a",
  1277 => x"e0c049bf",
  1278 => x"6a972966",
  1279 => x"9871484a",
  1280 => x"58a6f0c0",
  1281 => x"81c4496e",
  1282 => x"66dc4d69",
  1283 => x"a866d848",
  1284 => x"87c8c002",
  1285 => x"c048a6d8",
  1286 => x"87c5c078",
  1287 => x"c148a6d8",
  1288 => x"1e66d878",
  1289 => x"751ee0c0",
  1290 => x"d6deff49",
  1291 => x"7086c887",
  1292 => x"acb7c04c",
  1293 => x"87d4c106",
  1294 => x"e0c08574",
  1295 => x"75897449",
  1296 => x"c6d5c14b",
  1297 => x"f1fe714a",
  1298 => x"85c287de",
  1299 => x"4866e8c0",
  1300 => x"ecc080c1",
  1301 => x"ecc058a6",
  1302 => x"81c14966",
  1303 => x"c002a970",
  1304 => x"a6d887c8",
  1305 => x"c078c048",
  1306 => x"a6d887c5",
  1307 => x"d878c148",
  1308 => x"a4c21e66",
  1309 => x"48e0c049",
  1310 => x"49708871",
  1311 => x"ff49751e",
  1312 => x"c887c0dd",
  1313 => x"a8b7c086",
  1314 => x"87c0ff01",
  1315 => x"0266e8c0",
  1316 => x"6e87d1c0",
  1317 => x"c081c949",
  1318 => x"6e5166e8",
  1319 => x"d7c0c148",
  1320 => x"87ccc078",
  1321 => x"81c9496e",
  1322 => x"486e51c2",
  1323 => x"78cbc1c1",
  1324 => x"c6c07ec1",
  1325 => x"f6dbff87",
  1326 => x"6e4c7087",
  1327 => x"87f5c002",
  1328 => x"c84866c4",
  1329 => x"c004a866",
  1330 => x"66c487cb",
  1331 => x"c880c148",
  1332 => x"e0c058a6",
  1333 => x"4866c887",
  1334 => x"a6cc88c1",
  1335 => x"87d5c058",
  1336 => x"05acc6c1",
  1337 => x"cc87c8c0",
  1338 => x"80c14866",
  1339 => x"ff58a6d0",
  1340 => x"7087fcda",
  1341 => x"4866d04c",
  1342 => x"a6d480c1",
  1343 => x"029c7458",
  1344 => x"c487cbc0",
  1345 => x"c8c14866",
  1346 => x"f204a866",
  1347 => x"daff87ff",
  1348 => x"66c487d4",
  1349 => x"03a8c748",
  1350 => x"c287e5c0",
  1351 => x"c048d0dc",
  1352 => x"4966c478",
  1353 => x"c0c191cb",
  1354 => x"a1c48166",
  1355 => x"c04a6a4a",
  1356 => x"66c47952",
  1357 => x"c880c148",
  1358 => x"a8c758a6",
  1359 => x"87dbff04",
  1360 => x"e08ed0ff",
  1361 => x"203a87fb",
  1362 => x"1e731e00",
  1363 => x"029b4b71",
  1364 => x"dcc287c6",
  1365 => x"78c048cc",
  1366 => x"dcc21ec7",
  1367 => x"1e49bfcc",
  1368 => x"1ef2d8c1",
  1369 => x"bfc8dcc2",
  1370 => x"87f4ee49",
  1371 => x"dcc286cc",
  1372 => x"e949bfc8",
  1373 => x"9b7387f9",
  1374 => x"c187c802",
  1375 => x"c049f2d8",
  1376 => x"ff87cce5",
  1377 => x"1e87fedf",
  1378 => x"48dbcdc2",
  1379 => x"dac150c0",
  1380 => x"c049bfd5",
  1381 => x"c087c8f3",
  1382 => x"1e4f2648",
  1383 => x"c187e5c7",
  1384 => x"87e5fe49",
  1385 => x"87fdf3fe",
  1386 => x"cd029870",
  1387 => x"d8fbfe87",
  1388 => x"02987087",
  1389 => x"4ac187c4",
  1390 => x"4ac087c2",
  1391 => x"ce059a72",
  1392 => x"c11ec087",
  1393 => x"c049efd7",
  1394 => x"c487d2f0",
  1395 => x"c087fe86",
  1396 => x"c087f2f6",
  1397 => x"fad7c11e",
  1398 => x"c0f0c049",
  1399 => x"fe1ec087",
  1400 => x"497087e5",
  1401 => x"87f5efc0",
  1402 => x"f887d8c3",
  1403 => x"534f268e",
  1404 => x"61662044",
  1405 => x"64656c69",
  1406 => x"6f42002e",
  1407 => x"6e69746f",
  1408 => x"2e2e2e67",
  1409 => x"e7c01e00",
  1410 => x"87fa87e1",
  1411 => x"c21e4f26",
  1412 => x"c048ccdc",
  1413 => x"c8dcc278",
  1414 => x"fd78c048",
  1415 => x"87e587fd",
  1416 => x"4f2648c0",
  1417 => x"78452080",
  1418 => x"80007469",
  1419 => x"63614220",
  1420 => x"0fc7006b",
  1421 => x"27210000",
  1422 => x"00000000",
  1423 => x"000fc700",
  1424 => x"00273f00",
  1425 => x"00000000",
  1426 => x"00000fc7",
  1427 => x"0000275d",
  1428 => x"c7000000",
  1429 => x"7b00000f",
  1430 => x"00000027",
  1431 => x"0fc70000",
  1432 => x"27990000",
  1433 => x"00000000",
  1434 => x"000fc700",
  1435 => x"0027b700",
  1436 => x"00000000",
  1437 => x"00000fc7",
  1438 => x"000027d5",
  1439 => x"c7000000",
  1440 => x"0000000f",
  1441 => x"00000000",
  1442 => x"105c0000",
  1443 => x"00000000",
  1444 => x"00000000",
  1445 => x"00169900",
  1446 => x"4f4f4200",
  1447 => x"20202054",
  1448 => x"4d4f5220",
  1449 => x"616f4c00",
  1450 => x"2e2a2064",
  1451 => x"f0fe1e00",
  1452 => x"cd78c048",
  1453 => x"26097909",
  1454 => x"fe1e1e4f",
  1455 => x"487ebff0",
  1456 => x"1e4f2626",
  1457 => x"c148f0fe",
  1458 => x"1e4f2678",
  1459 => x"c048f0fe",
  1460 => x"1e4f2678",
  1461 => x"52c04a71",
  1462 => x"0e4f2652",
  1463 => x"5d5c5b5e",
  1464 => x"7186f40e",
  1465 => x"7e6d974d",
  1466 => x"974ca5c1",
  1467 => x"a6c8486c",
  1468 => x"c4486e58",
  1469 => x"c505a866",
  1470 => x"c048ff87",
  1471 => x"caff87e6",
  1472 => x"49a5c287",
  1473 => x"714b6c97",
  1474 => x"6b974ba3",
  1475 => x"7e6c974b",
  1476 => x"80c1486e",
  1477 => x"c758a6c8",
  1478 => x"58a6cc98",
  1479 => x"fe7c9770",
  1480 => x"487387e1",
  1481 => x"4d268ef4",
  1482 => x"4b264c26",
  1483 => x"5e0e4f26",
  1484 => x"f40e5c5b",
  1485 => x"d84c7186",
  1486 => x"ffc34a66",
  1487 => x"4ba4c29a",
  1488 => x"73496c97",
  1489 => x"517249a1",
  1490 => x"6e7e6c97",
  1491 => x"c880c148",
  1492 => x"98c758a6",
  1493 => x"7058a6cc",
  1494 => x"ff8ef454",
  1495 => x"1e1e87ca",
  1496 => x"e087e8fd",
  1497 => x"c0494abf",
  1498 => x"0299c0e0",
  1499 => x"1e7287cb",
  1500 => x"49f3dfc2",
  1501 => x"c487f7fe",
  1502 => x"87fdfc86",
  1503 => x"c2fd7e70",
  1504 => x"4f262687",
  1505 => x"f3dfc21e",
  1506 => x"87c7fd49",
  1507 => x"49deddc1",
  1508 => x"c587dafc",
  1509 => x"4f2687d9",
  1510 => x"5c5b5e0e",
  1511 => x"e0c20e5d",
  1512 => x"c14abfd2",
  1513 => x"49bfecdf",
  1514 => x"71bc724c",
  1515 => x"87dbfc4d",
  1516 => x"49744bc0",
  1517 => x"d50299d0",
  1518 => x"d0497587",
  1519 => x"c01e7199",
  1520 => x"fee5c11e",
  1521 => x"1282734a",
  1522 => x"87e4c049",
  1523 => x"2cc186c8",
  1524 => x"abc8832d",
  1525 => x"87daff04",
  1526 => x"c187e8fb",
  1527 => x"c248ecdf",
  1528 => x"78bfd2e0",
  1529 => x"4c264d26",
  1530 => x"4f264b26",
  1531 => x"00000000",
  1532 => x"48d0ff1e",
  1533 => x"ff78e1c8",
  1534 => x"78c548d4",
  1535 => x"c30266c4",
  1536 => x"78e0c387",
  1537 => x"c60266c8",
  1538 => x"48d4ff87",
  1539 => x"ff78f0c3",
  1540 => x"787148d4",
  1541 => x"c848d0ff",
  1542 => x"e0c078e1",
  1543 => x"0e4f2678",
  1544 => x"0e5c5b5e",
  1545 => x"dfc24c71",
  1546 => x"eefa49f3",
  1547 => x"c04a7087",
  1548 => x"c204aab7",
  1549 => x"e0c387e3",
  1550 => x"87c905aa",
  1551 => x"48e2e3c1",
  1552 => x"d4c278c1",
  1553 => x"aaf0c387",
  1554 => x"c187c905",
  1555 => x"c148dee3",
  1556 => x"87f5c178",
  1557 => x"bfe2e3c1",
  1558 => x"7287c702",
  1559 => x"b3c0c24b",
  1560 => x"4b7287c2",
  1561 => x"d1059c74",
  1562 => x"dee3c187",
  1563 => x"e3c11ebf",
  1564 => x"721ebfe2",
  1565 => x"87f8fd49",
  1566 => x"e3c186c8",
  1567 => x"c002bfde",
  1568 => x"497387e0",
  1569 => x"9129b7c4",
  1570 => x"81fee4c1",
  1571 => x"9acf4a73",
  1572 => x"48c192c2",
  1573 => x"4a703072",
  1574 => x"4872baff",
  1575 => x"79709869",
  1576 => x"497387db",
  1577 => x"9129b7c4",
  1578 => x"81fee4c1",
  1579 => x"9acf4a73",
  1580 => x"48c392c2",
  1581 => x"4a703072",
  1582 => x"70b06948",
  1583 => x"e2e3c179",
  1584 => x"c178c048",
  1585 => x"c048dee3",
  1586 => x"f3dfc278",
  1587 => x"87cbf849",
  1588 => x"b7c04a70",
  1589 => x"ddfd03aa",
  1590 => x"fc48c087",
  1591 => x"000087c8",
  1592 => x"00000000",
  1593 => x"711e0000",
  1594 => x"f2fc494a",
  1595 => x"1e4f2687",
  1596 => x"49724ac0",
  1597 => x"e4c191c4",
  1598 => x"79c081fe",
  1599 => x"b7d082c1",
  1600 => x"87ee04aa",
  1601 => x"5e0e4f26",
  1602 => x"0e5d5c5b",
  1603 => x"faf64d71",
  1604 => x"c44a7587",
  1605 => x"c1922ab7",
  1606 => x"7582fee4",
  1607 => x"c29ccf4c",
  1608 => x"4b496a94",
  1609 => x"9bc32b74",
  1610 => x"307448c2",
  1611 => x"bcff4c70",
  1612 => x"98714874",
  1613 => x"caf67a70",
  1614 => x"fa487387",
  1615 => x"000087e6",
  1616 => x"00000000",
  1617 => x"00000000",
  1618 => x"00000000",
  1619 => x"00000000",
  1620 => x"00000000",
  1621 => x"00000000",
  1622 => x"00000000",
  1623 => x"00000000",
  1624 => x"00000000",
  1625 => x"00000000",
  1626 => x"00000000",
  1627 => x"00000000",
  1628 => x"00000000",
  1629 => x"00000000",
  1630 => x"00000000",
  1631 => x"1e160000",
  1632 => x"362e2526",
  1633 => x"ff1e3e3d",
  1634 => x"e1c848d0",
  1635 => x"ff487178",
  1636 => x"c47808d4",
  1637 => x"d4ff4866",
  1638 => x"4f267808",
  1639 => x"c44a711e",
  1640 => x"e0c11e66",
  1641 => x"ddff49a2",
  1642 => x"4966c887",
  1643 => x"ff29b7c8",
  1644 => x"787148d4",
  1645 => x"c048d0ff",
  1646 => x"262678e0",
  1647 => x"d4ff1e4f",
  1648 => x"7affc34a",
  1649 => x"c848d0ff",
  1650 => x"7ade78e1",
  1651 => x"bffddfc2",
  1652 => x"c848497a",
  1653 => x"717a7028",
  1654 => x"7028d048",
  1655 => x"d848717a",
  1656 => x"ff7a7028",
  1657 => x"e0c048d0",
  1658 => x"0e4f2678",
  1659 => x"5d5c5b5e",
  1660 => x"c24c710e",
  1661 => x"4dbffddf",
  1662 => x"d02b744b",
  1663 => x"83c19b66",
  1664 => x"04ab66d4",
  1665 => x"4bc087c2",
  1666 => x"66d04a74",
  1667 => x"ff317249",
  1668 => x"739975b9",
  1669 => x"70307248",
  1670 => x"b071484a",
  1671 => x"58c1e0c2",
  1672 => x"2687dafe",
  1673 => x"264c264d",
  1674 => x"1e4f264b",
  1675 => x"c848d0ff",
  1676 => x"487178c9",
  1677 => x"7808d4ff",
  1678 => x"711e4f26",
  1679 => x"87eb494a",
  1680 => x"c848d0ff",
  1681 => x"1e4f2678",
  1682 => x"4b711e73",
  1683 => x"bfcde0c2",
  1684 => x"c287c302",
  1685 => x"d0ff87eb",
  1686 => x"78c9c848",
  1687 => x"e0c04973",
  1688 => x"48d4ffb1",
  1689 => x"e0c27871",
  1690 => x"78c048c1",
  1691 => x"c50266c8",
  1692 => x"49ffc387",
  1693 => x"49c087c2",
  1694 => x"59c9e0c2",
  1695 => x"c60266cc",
  1696 => x"d5d5c587",
  1697 => x"cf87c44a",
  1698 => x"c24affff",
  1699 => x"c25acde0",
  1700 => x"c148cde0",
  1701 => x"2687c478",
  1702 => x"264c264d",
  1703 => x"0e4f264b",
  1704 => x"5d5c5b5e",
  1705 => x"c24a710e",
  1706 => x"4cbfc9e0",
  1707 => x"cb029a72",
  1708 => x"91c84987",
  1709 => x"4bfde8c1",
  1710 => x"87c48371",
  1711 => x"4bfdecc1",
  1712 => x"49134dc0",
  1713 => x"e0c29974",
  1714 => x"ffb9bfc5",
  1715 => x"787148d4",
  1716 => x"852cb7c1",
  1717 => x"04adb7c8",
  1718 => x"e0c287e8",
  1719 => x"c848bfc1",
  1720 => x"c5e0c280",
  1721 => x"87effe58",
  1722 => x"711e731e",
  1723 => x"9a4a134b",
  1724 => x"7287cb02",
  1725 => x"87e7fe49",
  1726 => x"059a4a13",
  1727 => x"dafe87f5",
  1728 => x"e0c21e87",
  1729 => x"c249bfc1",
  1730 => x"c148c1e0",
  1731 => x"c0c478a1",
  1732 => x"db03a9b7",
  1733 => x"48d4ff87",
  1734 => x"bfc5e0c2",
  1735 => x"c1e0c278",
  1736 => x"e0c249bf",
  1737 => x"a1c148c1",
  1738 => x"b7c0c478",
  1739 => x"87e504a9",
  1740 => x"c848d0ff",
  1741 => x"cde0c278",
  1742 => x"2678c048",
  1743 => x"0000004f",
  1744 => x"00000000",
  1745 => x"00000000",
  1746 => x"00005f5f",
  1747 => x"03030000",
  1748 => x"00030300",
  1749 => x"7f7f1400",
  1750 => x"147f7f14",
  1751 => x"2e240000",
  1752 => x"123a6b6b",
  1753 => x"366a4c00",
  1754 => x"32566c18",
  1755 => x"4f7e3000",
  1756 => x"683a7759",
  1757 => x"04000040",
  1758 => x"00000307",
  1759 => x"1c000000",
  1760 => x"0041633e",
  1761 => x"41000000",
  1762 => x"001c3e63",
  1763 => x"3e2a0800",
  1764 => x"2a3e1c1c",
  1765 => x"08080008",
  1766 => x"08083e3e",
  1767 => x"80000000",
  1768 => x"000060e0",
  1769 => x"08080000",
  1770 => x"08080808",
  1771 => x"00000000",
  1772 => x"00006060",
  1773 => x"30604000",
  1774 => x"03060c18",
  1775 => x"7f3e0001",
  1776 => x"3e7f4d59",
  1777 => x"06040000",
  1778 => x"00007f7f",
  1779 => x"63420000",
  1780 => x"464f5971",
  1781 => x"63220000",
  1782 => x"367f4949",
  1783 => x"161c1800",
  1784 => x"107f7f13",
  1785 => x"67270000",
  1786 => x"397d4545",
  1787 => x"7e3c0000",
  1788 => x"3079494b",
  1789 => x"01010000",
  1790 => x"070f7971",
  1791 => x"7f360000",
  1792 => x"367f4949",
  1793 => x"4f060000",
  1794 => x"1e3f6949",
  1795 => x"00000000",
  1796 => x"00006666",
  1797 => x"80000000",
  1798 => x"000066e6",
  1799 => x"08080000",
  1800 => x"22221414",
  1801 => x"14140000",
  1802 => x"14141414",
  1803 => x"22220000",
  1804 => x"08081414",
  1805 => x"03020000",
  1806 => x"060f5951",
  1807 => x"417f3e00",
  1808 => x"1e1f555d",
  1809 => x"7f7e0000",
  1810 => x"7e7f0909",
  1811 => x"7f7f0000",
  1812 => x"367f4949",
  1813 => x"3e1c0000",
  1814 => x"41414163",
  1815 => x"7f7f0000",
  1816 => x"1c3e6341",
  1817 => x"7f7f0000",
  1818 => x"41414949",
  1819 => x"7f7f0000",
  1820 => x"01010909",
  1821 => x"7f3e0000",
  1822 => x"7a7b4941",
  1823 => x"7f7f0000",
  1824 => x"7f7f0808",
  1825 => x"41000000",
  1826 => x"00417f7f",
  1827 => x"60200000",
  1828 => x"3f7f4040",
  1829 => x"087f7f00",
  1830 => x"4163361c",
  1831 => x"7f7f0000",
  1832 => x"40404040",
  1833 => x"067f7f00",
  1834 => x"7f7f060c",
  1835 => x"067f7f00",
  1836 => x"7f7f180c",
  1837 => x"7f3e0000",
  1838 => x"3e7f4141",
  1839 => x"7f7f0000",
  1840 => x"060f0909",
  1841 => x"417f3e00",
  1842 => x"407e7f61",
  1843 => x"7f7f0000",
  1844 => x"667f1909",
  1845 => x"6f260000",
  1846 => x"327b594d",
  1847 => x"01010000",
  1848 => x"01017f7f",
  1849 => x"7f3f0000",
  1850 => x"3f7f4040",
  1851 => x"3f0f0000",
  1852 => x"0f3f7070",
  1853 => x"307f7f00",
  1854 => x"7f7f3018",
  1855 => x"36634100",
  1856 => x"63361c1c",
  1857 => x"06030141",
  1858 => x"03067c7c",
  1859 => x"59716101",
  1860 => x"4143474d",
  1861 => x"7f000000",
  1862 => x"0041417f",
  1863 => x"06030100",
  1864 => x"6030180c",
  1865 => x"41000040",
  1866 => x"007f7f41",
  1867 => x"060c0800",
  1868 => x"080c0603",
  1869 => x"80808000",
  1870 => x"80808080",
  1871 => x"00000000",
  1872 => x"00040703",
  1873 => x"74200000",
  1874 => x"787c5454",
  1875 => x"7f7f0000",
  1876 => x"387c4444",
  1877 => x"7c380000",
  1878 => x"00444444",
  1879 => x"7c380000",
  1880 => x"7f7f4444",
  1881 => x"7c380000",
  1882 => x"185c5454",
  1883 => x"7e040000",
  1884 => x"0005057f",
  1885 => x"bc180000",
  1886 => x"7cfca4a4",
  1887 => x"7f7f0000",
  1888 => x"787c0404",
  1889 => x"00000000",
  1890 => x"00407d3d",
  1891 => x"80800000",
  1892 => x"007dfd80",
  1893 => x"7f7f0000",
  1894 => x"446c3810",
  1895 => x"00000000",
  1896 => x"00407f3f",
  1897 => x"0c7c7c00",
  1898 => x"787c0c18",
  1899 => x"7c7c0000",
  1900 => x"787c0404",
  1901 => x"7c380000",
  1902 => x"387c4444",
  1903 => x"fcfc0000",
  1904 => x"183c2424",
  1905 => x"3c180000",
  1906 => x"fcfc2424",
  1907 => x"7c7c0000",
  1908 => x"080c0404",
  1909 => x"5c480000",
  1910 => x"20745454",
  1911 => x"3f040000",
  1912 => x"0044447f",
  1913 => x"7c3c0000",
  1914 => x"7c7c4040",
  1915 => x"3c1c0000",
  1916 => x"1c3c6060",
  1917 => x"607c3c00",
  1918 => x"3c7c6030",
  1919 => x"386c4400",
  1920 => x"446c3810",
  1921 => x"bc1c0000",
  1922 => x"1c3c60e0",
  1923 => x"64440000",
  1924 => x"444c5c74",
  1925 => x"08080000",
  1926 => x"4141773e",
  1927 => x"00000000",
  1928 => x"00007f7f",
  1929 => x"41410000",
  1930 => x"08083e77",
  1931 => x"01010200",
  1932 => x"01020203",
  1933 => x"7f7f7f00",
  1934 => x"7f7f7f7f",
  1935 => x"1c080800",
  1936 => x"7f3e3e1c",
  1937 => x"3e7f7f7f",
  1938 => x"081c1c3e",
  1939 => x"18100008",
  1940 => x"10187c7c",
  1941 => x"30100000",
  1942 => x"10307c7c",
  1943 => x"60301000",
  1944 => x"061e7860",
  1945 => x"3c664200",
  1946 => x"42663c18",
  1947 => x"6a387800",
  1948 => x"386cc6c2",
  1949 => x"00006000",
  1950 => x"60000060",
  1951 => x"5b5e0e00",
  1952 => x"1e0e5d5c",
  1953 => x"e0c24c71",
  1954 => x"c04dbfde",
  1955 => x"741ec04b",
  1956 => x"87c702ab",
  1957 => x"c048a6c4",
  1958 => x"c487c578",
  1959 => x"78c148a6",
  1960 => x"731e66c4",
  1961 => x"87dfee49",
  1962 => x"e0c086c8",
  1963 => x"87efef49",
  1964 => x"6a4aa5c4",
  1965 => x"87f0f049",
  1966 => x"cb87c6f1",
  1967 => x"c883c185",
  1968 => x"ff04abb7",
  1969 => x"262687c7",
  1970 => x"264c264d",
  1971 => x"1e4f264b",
  1972 => x"e0c24a71",
  1973 => x"e0c25ae2",
  1974 => x"78c748e2",
  1975 => x"87ddfe49",
  1976 => x"731e4f26",
  1977 => x"c04a711e",
  1978 => x"d303aab7",
  1979 => x"f2c8c287",
  1980 => x"87c405bf",
  1981 => x"87c24bc1",
  1982 => x"c8c24bc0",
  1983 => x"87c45bf6",
  1984 => x"5af6c8c2",
  1985 => x"bff2c8c2",
  1986 => x"c19ac14a",
  1987 => x"ec49a2c0",
  1988 => x"48fc87e8",
  1989 => x"bff2c8c2",
  1990 => x"87effe78",
  1991 => x"c44a711e",
  1992 => x"49721e66",
  1993 => x"2687f5e9",
  1994 => x"c21e4f26",
  1995 => x"49bff2c8",
  1996 => x"c287f3e6",
  1997 => x"e848d6e0",
  1998 => x"e0c278bf",
  1999 => x"bfec48d2",
  2000 => x"d6e0c278",
  2001 => x"c3494abf",
  2002 => x"b7c899ff",
  2003 => x"7148722a",
  2004 => x"dee0c2b0",
  2005 => x"0e4f2658",
  2006 => x"5d5c5b5e",
  2007 => x"ff4b710e",
  2008 => x"e0c287c8",
  2009 => x"50c048d1",
  2010 => x"d9e64973",
  2011 => x"4c497087",
  2012 => x"eecb9cc2",
  2013 => x"87c2cb49",
  2014 => x"c24d4970",
  2015 => x"bf97d1e0",
  2016 => x"87e2c105",
  2017 => x"c24966d0",
  2018 => x"99bfdae0",
  2019 => x"d487d605",
  2020 => x"e0c24966",
  2021 => x"0599bfd2",
  2022 => x"497387cb",
  2023 => x"7087e7e5",
  2024 => x"c1c10298",
  2025 => x"fe4cc187",
  2026 => x"497587c0",
  2027 => x"7087d7ca",
  2028 => x"87c60298",
  2029 => x"48d1e0c2",
  2030 => x"e0c250c1",
  2031 => x"05bf97d1",
  2032 => x"c287e3c0",
  2033 => x"49bfdae0",
  2034 => x"059966d0",
  2035 => x"c287d6ff",
  2036 => x"49bfd2e0",
  2037 => x"059966d4",
  2038 => x"7387caff",
  2039 => x"87e6e449",
  2040 => x"fe059870",
  2041 => x"487487ff",
  2042 => x"0e87dcfb",
  2043 => x"5d5c5b5e",
  2044 => x"c086f40e",
  2045 => x"bfec4c4d",
  2046 => x"48a6c47e",
  2047 => x"bfdee0c2",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
